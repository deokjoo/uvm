
//
//
//
//
//

class axis_agent_cfg extends uvm_object;
    `uvm_object_utils(axis_agent_cfg)

    function new(string name="axis_agent_cfg");
        super.new(name);
    endfunction

endclass



