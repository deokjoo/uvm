//
//
//
//
//
//


package axis_test_pkg;
    `include "uvm_macros.svh"
    
    import uvm_pkg::*;


    // test class
    `include "axis_base_test.svh"

endpackage