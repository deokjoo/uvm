//
//
//
//
//

class filter_env_cfg extends uvm_object;
    `uvm_object_utils(filter_env_cfg)

    function new(string name="filter_env_cfg");
        super.new(name);
    endfunction

endclass

//
//

