//
//
//
//
//

class axis_agent extends uvm_agent;
    `uvm_component_utils(axis_agent)

    function new (string name="axis_agent", uvm_component parent=null);
        super.new(name, parent);
    endfunction

endclass

//
//
