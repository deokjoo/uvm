//
//
//
//
//
//

class axis_base_test extends uvm_test;
    `uvm_component_utils(axis_base_test)

    //        
    // constructor
    function new(string name="axis_base_test", uvm_component parent=null);
       super.new(name, parent);    
    endfunction

    //


endclass
