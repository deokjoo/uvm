//
//
//
//
//
//
package axis_test_pkg;
    `include "uvm_macros.svh"
    
    import uvm_pkg::*;

    //agent

    `include "axis_agent.svh"
    // env
    `include "filter_env_cfg.svh"
    `include "filter_env.svh"

    //test
    `include "axis_base_test.svh"

endpackage


